// soc_system.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        clk_clk,                               //          clk.clk
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK, // hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,   //             .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,   //             .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,   //             .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,   //             .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,   //             .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,   //             .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,    //             .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL, //             .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL, //             .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK, //             .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,   //             .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,   //             .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,   //             .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,     //             .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,     //             .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,     //             .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,     //             .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,     //             .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,     //             .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,     //             .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,      //             .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,      //             .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,     //             .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,      //             .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,      //             .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,      //             .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,      //             .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,      //             .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,      //             .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,      //             .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,      //             .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,      //             .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,      //             .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,     //             .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,     //             .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,     //             .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,     //             .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim0_inst_CLK,    //             .hps_io_spim0_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim0_inst_MOSI,   //             .hps_io_spim0_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim0_inst_MISO,   //             .hps_io_spim0_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim0_inst_SS0,    //             .hps_io_spim0_inst_SS0
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,    //             .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,   //             .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,   //             .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,    //             .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,     //             .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,     //             .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,     //             .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,     //             .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,     //             .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,     //             .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,  //             .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,  //             .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO37,  //             .hps_io_gpio_inst_GPIO37
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,  //             .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,  //             .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO44,  //             .hps_io_gpio_inst_GPIO44
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,  //             .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,  //             .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,  //             .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,  //             .hps_io_gpio_inst_GPIO61
		output wire [14:0] memory_mem_a,                          //       memory.mem_a
		output wire [2:0]  memory_mem_ba,                         //             .mem_ba
		output wire        memory_mem_ck,                         //             .mem_ck
		output wire        memory_mem_ck_n,                       //             .mem_ck_n
		output wire        memory_mem_cke,                        //             .mem_cke
		output wire        memory_mem_cs_n,                       //             .mem_cs_n
		output wire        memory_mem_ras_n,                      //             .mem_ras_n
		output wire        memory_mem_cas_n,                      //             .mem_cas_n
		output wire        memory_mem_we_n,                       //             .mem_we_n
		output wire        memory_mem_reset_n,                    //             .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                         //             .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                        //             .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                      //             .mem_dqs_n
		output wire        memory_mem_odt,                        //             .mem_odt
		output wire [3:0]  memory_mem_dm,                         //             .mem_dm
		input  wire        memory_oct_rzqin,                      //             .oct_rzqin
		input  wire [31:0] pp_in_axi_export,                      //    pp_in_axi.export
		output wire [31:0] pp_out_axi_export                      //   pp_out_axi.export
	);

	wire          hps_0_h2f_reset_reset;                                                         // hps_0:h2f_rst_n -> rst_controller:reset_in0
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                                  // hps_0:h2f_AWBURST -> mm_interconnect_0:hps_0_h2f_axi_master_awburst
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                                    // hps_0:h2f_ARLEN -> mm_interconnect_0:hps_0_h2f_axi_master_arlen
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                                    // hps_0:h2f_WSTRB -> mm_interconnect_0:hps_0_h2f_axi_master_wstrb
	wire          hps_0_h2f_axi_master_wready;                                                   // mm_interconnect_0:hps_0_h2f_axi_master_wready -> hps_0:h2f_WREADY
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                      // mm_interconnect_0:hps_0_h2f_axi_master_rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_rready;                                                   // hps_0:h2f_RREADY -> mm_interconnect_0:hps_0_h2f_axi_master_rready
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                                    // hps_0:h2f_AWLEN -> mm_interconnect_0:hps_0_h2f_axi_master_awlen
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                      // hps_0:h2f_WID -> mm_interconnect_0:hps_0_h2f_axi_master_wid
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                                  // hps_0:h2f_ARCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_arcache
	wire          hps_0_h2f_axi_master_wvalid;                                                   // hps_0:h2f_WVALID -> mm_interconnect_0:hps_0_h2f_axi_master_wvalid
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                                   // hps_0:h2f_ARADDR -> mm_interconnect_0:hps_0_h2f_axi_master_araddr
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                                   // hps_0:h2f_ARPROT -> mm_interconnect_0:hps_0_h2f_axi_master_arprot
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                                   // hps_0:h2f_AWPROT -> mm_interconnect_0:hps_0_h2f_axi_master_awprot
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                                    // hps_0:h2f_WDATA -> mm_interconnect_0:hps_0_h2f_axi_master_wdata
	wire          hps_0_h2f_axi_master_arvalid;                                                  // hps_0:h2f_ARVALID -> mm_interconnect_0:hps_0_h2f_axi_master_arvalid
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                                  // hps_0:h2f_AWCACHE -> mm_interconnect_0:hps_0_h2f_axi_master_awcache
	wire   [11:0] hps_0_h2f_axi_master_arid;                                                     // hps_0:h2f_ARID -> mm_interconnect_0:hps_0_h2f_axi_master_arid
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                                   // hps_0:h2f_ARLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_arlock
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                                   // hps_0:h2f_AWLOCK -> mm_interconnect_0:hps_0_h2f_axi_master_awlock
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                                   // hps_0:h2f_AWADDR -> mm_interconnect_0:hps_0_h2f_axi_master_awaddr
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                                    // mm_interconnect_0:hps_0_h2f_axi_master_bresp -> hps_0:h2f_BRESP
	wire          hps_0_h2f_axi_master_arready;                                                  // mm_interconnect_0:hps_0_h2f_axi_master_arready -> hps_0:h2f_ARREADY
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                                    // mm_interconnect_0:hps_0_h2f_axi_master_rdata -> hps_0:h2f_RDATA
	wire          hps_0_h2f_axi_master_awready;                                                  // mm_interconnect_0:hps_0_h2f_axi_master_awready -> hps_0:h2f_AWREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                                  // hps_0:h2f_ARBURST -> mm_interconnect_0:hps_0_h2f_axi_master_arburst
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                                   // hps_0:h2f_ARSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_arsize
	wire          hps_0_h2f_axi_master_bready;                                                   // hps_0:h2f_BREADY -> mm_interconnect_0:hps_0_h2f_axi_master_bready
	wire          hps_0_h2f_axi_master_rlast;                                                    // mm_interconnect_0:hps_0_h2f_axi_master_rlast -> hps_0:h2f_RLAST
	wire          hps_0_h2f_axi_master_wlast;                                                    // hps_0:h2f_WLAST -> mm_interconnect_0:hps_0_h2f_axi_master_wlast
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                                    // mm_interconnect_0:hps_0_h2f_axi_master_rresp -> hps_0:h2f_RRESP
	wire   [11:0] hps_0_h2f_axi_master_awid;                                                     // hps_0:h2f_AWID -> mm_interconnect_0:hps_0_h2f_axi_master_awid
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                      // mm_interconnect_0:hps_0_h2f_axi_master_bid -> hps_0:h2f_BID
	wire          hps_0_h2f_axi_master_bvalid;                                                   // mm_interconnect_0:hps_0_h2f_axi_master_bvalid -> hps_0:h2f_BVALID
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                                   // hps_0:h2f_AWSIZE -> mm_interconnect_0:hps_0_h2f_axi_master_awsize
	wire          hps_0_h2f_axi_master_awvalid;                                                  // hps_0:h2f_AWVALID -> mm_interconnect_0:hps_0_h2f_axi_master_awvalid
	wire          hps_0_h2f_axi_master_rvalid;                                                   // mm_interconnect_0:hps_0_h2f_axi_master_rvalid -> hps_0:h2f_RVALID
	wire          mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_chipselect; // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_chipselect -> parallel_port_out_axi:chipselect
	wire   [31:0] mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_readdata;   // parallel_port_out_axi:readdata -> mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_readdata
	wire    [1:0] mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_address;    // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_address -> parallel_port_out_axi:address
	wire          mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_read;       // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_read -> parallel_port_out_axi:read
	wire    [3:0] mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_byteenable; // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_byteenable -> parallel_port_out_axi:byteenable
	wire          mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_write;      // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_write -> parallel_port_out_axi:write
	wire   [31:0] mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_writedata;  // mm_interconnect_0:parallel_port_out_axi_avalon_parallel_port_slave_writedata -> parallel_port_out_axi:writedata
	wire          mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_chipselect;  // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_chipselect -> parallel_port_in_axi:chipselect
	wire   [31:0] mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_readdata;    // parallel_port_in_axi:readdata -> mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_readdata
	wire    [1:0] mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_address;     // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_address -> parallel_port_in_axi:address
	wire          mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_read;        // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_read -> parallel_port_in_axi:read
	wire    [3:0] mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_byteenable;  // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_byteenable -> parallel_port_in_axi:byteenable
	wire          mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_write;       // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_write -> parallel_port_in_axi:write
	wire   [31:0] mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_writedata;   // mm_interconnect_0:parallel_port_in_axi_avalon_parallel_port_slave_writedata -> parallel_port_in_axi:writedata
	wire   [31:0] hps_0_f2h_irq0_irq;                                                            // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                            // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                                // rst_controller:reset_out -> [mm_interconnect_0:parallel_port_out_axi_reset_reset_bridge_in_reset_reset, parallel_port_in_axi:reset, parallel_port_out_axi:reset]

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                          //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                         //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                         //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                       //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                        //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                       //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                      //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                      //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                       //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                    //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                         //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                        //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                      //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                        //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                         //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                      //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK), //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL), //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL), //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK), //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),     //                  .hps_io_usb1_inst_NXT
		.hps_io_spim0_inst_CLK    (hps_0_hps_io_hps_io_spim0_inst_CLK),    //                  .hps_io_spim0_inst_CLK
		.hps_io_spim0_inst_MOSI   (hps_0_hps_io_hps_io_spim0_inst_MOSI),   //                  .hps_io_spim0_inst_MOSI
		.hps_io_spim0_inst_MISO   (hps_0_hps_io_hps_io_spim0_inst_MISO),   //                  .hps_io_spim0_inst_MISO
		.hps_io_spim0_inst_SS0    (hps_0_hps_io_hps_io_spim0_inst_SS0),    //                  .hps_io_spim0_inst_SS0
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),    //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),   //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),   //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),    //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO37  (hps_0_hps_io_hps_io_gpio_inst_GPIO37),  //                  .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),  //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO44  (hps_0_hps_io_hps_io_gpio_inst_GPIO44),  //                  .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),  //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),                 //         h2f_reset.reset_n
		.f2h_sdram0_clk           (clk_clk),                               //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (),                                      //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (),                                      //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (),                                      //                  .waitrequest
		.f2h_sdram0_READDATA      (),                                      //                  .readdata
		.f2h_sdram0_READDATAVALID (),                                      //                  .readdatavalid
		.f2h_sdram0_READ          (),                                      //                  .read
		.f2h_sdram0_WRITEDATA     (),                                      //                  .writedata
		.f2h_sdram0_BYTEENABLE    (),                                      //                  .byteenable
		.f2h_sdram0_WRITE         (),                                      //                  .write
		.h2f_axi_clk              (clk_clk),                               //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),             //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),           //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),            //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),           //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),          //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),           //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),          //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),           //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),          //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),          //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),              //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),            //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),            //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),            //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),           //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),           //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),              //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),            //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),           //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),           //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),             //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),           //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),            //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),           //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),          //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),           //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),          //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),           //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),          //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),          //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),              //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),            //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),            //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),            //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),           //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),           //                  .rready
		.f2h_axi_clk              (clk_clk),                               //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                      //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                      //                  .awaddr
		.f2h_AWLEN                (),                                      //                  .awlen
		.f2h_AWSIZE               (),                                      //                  .awsize
		.f2h_AWBURST              (),                                      //                  .awburst
		.f2h_AWLOCK               (),                                      //                  .awlock
		.f2h_AWCACHE              (),                                      //                  .awcache
		.f2h_AWPROT               (),                                      //                  .awprot
		.f2h_AWVALID              (),                                      //                  .awvalid
		.f2h_AWREADY              (),                                      //                  .awready
		.f2h_AWUSER               (),                                      //                  .awuser
		.f2h_WID                  (),                                      //                  .wid
		.f2h_WDATA                (),                                      //                  .wdata
		.f2h_WSTRB                (),                                      //                  .wstrb
		.f2h_WLAST                (),                                      //                  .wlast
		.f2h_WVALID               (),                                      //                  .wvalid
		.f2h_WREADY               (),                                      //                  .wready
		.f2h_BID                  (),                                      //                  .bid
		.f2h_BRESP                (),                                      //                  .bresp
		.f2h_BVALID               (),                                      //                  .bvalid
		.f2h_BREADY               (),                                      //                  .bready
		.f2h_ARID                 (),                                      //                  .arid
		.f2h_ARADDR               (),                                      //                  .araddr
		.f2h_ARLEN                (),                                      //                  .arlen
		.f2h_ARSIZE               (),                                      //                  .arsize
		.f2h_ARBURST              (),                                      //                  .arburst
		.f2h_ARLOCK               (),                                      //                  .arlock
		.f2h_ARCACHE              (),                                      //                  .arcache
		.f2h_ARPROT               (),                                      //                  .arprot
		.f2h_ARVALID              (),                                      //                  .arvalid
		.f2h_ARREADY              (),                                      //                  .arready
		.f2h_ARUSER               (),                                      //                  .aruser
		.f2h_RID                  (),                                      //                  .rid
		.f2h_RDATA                (),                                      //                  .rdata
		.f2h_RRESP                (),                                      //                  .rresp
		.f2h_RLAST                (),                                      //                  .rlast
		.f2h_RVALID               (),                                      //                  .rvalid
		.f2h_RREADY               (),                                      //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                               //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (),                                      // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (),                                      //                  .awaddr
		.h2f_lw_AWLEN             (),                                      //                  .awlen
		.h2f_lw_AWSIZE            (),                                      //                  .awsize
		.h2f_lw_AWBURST           (),                                      //                  .awburst
		.h2f_lw_AWLOCK            (),                                      //                  .awlock
		.h2f_lw_AWCACHE           (),                                      //                  .awcache
		.h2f_lw_AWPROT            (),                                      //                  .awprot
		.h2f_lw_AWVALID           (),                                      //                  .awvalid
		.h2f_lw_AWREADY           (),                                      //                  .awready
		.h2f_lw_WID               (),                                      //                  .wid
		.h2f_lw_WDATA             (),                                      //                  .wdata
		.h2f_lw_WSTRB             (),                                      //                  .wstrb
		.h2f_lw_WLAST             (),                                      //                  .wlast
		.h2f_lw_WVALID            (),                                      //                  .wvalid
		.h2f_lw_WREADY            (),                                      //                  .wready
		.h2f_lw_BID               (),                                      //                  .bid
		.h2f_lw_BRESP             (),                                      //                  .bresp
		.h2f_lw_BVALID            (),                                      //                  .bvalid
		.h2f_lw_BREADY            (),                                      //                  .bready
		.h2f_lw_ARID              (),                                      //                  .arid
		.h2f_lw_ARADDR            (),                                      //                  .araddr
		.h2f_lw_ARLEN             (),                                      //                  .arlen
		.h2f_lw_ARSIZE            (),                                      //                  .arsize
		.h2f_lw_ARBURST           (),                                      //                  .arburst
		.h2f_lw_ARLOCK            (),                                      //                  .arlock
		.h2f_lw_ARCACHE           (),                                      //                  .arcache
		.h2f_lw_ARPROT            (),                                      //                  .arprot
		.h2f_lw_ARVALID           (),                                      //                  .arvalid
		.h2f_lw_ARREADY           (),                                      //                  .arready
		.h2f_lw_RID               (),                                      //                  .rid
		.h2f_lw_RDATA             (),                                      //                  .rdata
		.h2f_lw_RRESP             (),                                      //                  .rresp
		.h2f_lw_RLAST             (),                                      //                  .rlast
		.h2f_lw_RVALID            (),                                      //                  .rvalid
		.h2f_lw_RREADY            (),                                      //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                    //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                     //          f2h_irq1.irq
	);

	soc_system_parallel_port_in_axi parallel_port_in_axi (
		.clk        (clk_clk),                                                                      //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                               //                      reset.reset
		.address    (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_readdata),   //                           .readdata
		.in_port    (pp_in_axi_export)                                                              //         external_interface.export
	);

	soc_system_parallel_port_out_axi parallel_port_out_axi (
		.clk        (clk_clk),                                                                       //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                                //                      reset.reset
		.address    (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_readdata),   //                           .readdata
		.out_port   (pp_out_axi_export)                                                              //         external_interface.export
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_axi_master_awid                                   (hps_0_h2f_axi_master_awid),                                                     //                              hps_0_h2f_axi_master.awid
		.hps_0_h2f_axi_master_awaddr                                 (hps_0_h2f_axi_master_awaddr),                                                   //                                                  .awaddr
		.hps_0_h2f_axi_master_awlen                                  (hps_0_h2f_axi_master_awlen),                                                    //                                                  .awlen
		.hps_0_h2f_axi_master_awsize                                 (hps_0_h2f_axi_master_awsize),                                                   //                                                  .awsize
		.hps_0_h2f_axi_master_awburst                                (hps_0_h2f_axi_master_awburst),                                                  //                                                  .awburst
		.hps_0_h2f_axi_master_awlock                                 (hps_0_h2f_axi_master_awlock),                                                   //                                                  .awlock
		.hps_0_h2f_axi_master_awcache                                (hps_0_h2f_axi_master_awcache),                                                  //                                                  .awcache
		.hps_0_h2f_axi_master_awprot                                 (hps_0_h2f_axi_master_awprot),                                                   //                                                  .awprot
		.hps_0_h2f_axi_master_awvalid                                (hps_0_h2f_axi_master_awvalid),                                                  //                                                  .awvalid
		.hps_0_h2f_axi_master_awready                                (hps_0_h2f_axi_master_awready),                                                  //                                                  .awready
		.hps_0_h2f_axi_master_wid                                    (hps_0_h2f_axi_master_wid),                                                      //                                                  .wid
		.hps_0_h2f_axi_master_wdata                                  (hps_0_h2f_axi_master_wdata),                                                    //                                                  .wdata
		.hps_0_h2f_axi_master_wstrb                                  (hps_0_h2f_axi_master_wstrb),                                                    //                                                  .wstrb
		.hps_0_h2f_axi_master_wlast                                  (hps_0_h2f_axi_master_wlast),                                                    //                                                  .wlast
		.hps_0_h2f_axi_master_wvalid                                 (hps_0_h2f_axi_master_wvalid),                                                   //                                                  .wvalid
		.hps_0_h2f_axi_master_wready                                 (hps_0_h2f_axi_master_wready),                                                   //                                                  .wready
		.hps_0_h2f_axi_master_bid                                    (hps_0_h2f_axi_master_bid),                                                      //                                                  .bid
		.hps_0_h2f_axi_master_bresp                                  (hps_0_h2f_axi_master_bresp),                                                    //                                                  .bresp
		.hps_0_h2f_axi_master_bvalid                                 (hps_0_h2f_axi_master_bvalid),                                                   //                                                  .bvalid
		.hps_0_h2f_axi_master_bready                                 (hps_0_h2f_axi_master_bready),                                                   //                                                  .bready
		.hps_0_h2f_axi_master_arid                                   (hps_0_h2f_axi_master_arid),                                                     //                                                  .arid
		.hps_0_h2f_axi_master_araddr                                 (hps_0_h2f_axi_master_araddr),                                                   //                                                  .araddr
		.hps_0_h2f_axi_master_arlen                                  (hps_0_h2f_axi_master_arlen),                                                    //                                                  .arlen
		.hps_0_h2f_axi_master_arsize                                 (hps_0_h2f_axi_master_arsize),                                                   //                                                  .arsize
		.hps_0_h2f_axi_master_arburst                                (hps_0_h2f_axi_master_arburst),                                                  //                                                  .arburst
		.hps_0_h2f_axi_master_arlock                                 (hps_0_h2f_axi_master_arlock),                                                   //                                                  .arlock
		.hps_0_h2f_axi_master_arcache                                (hps_0_h2f_axi_master_arcache),                                                  //                                                  .arcache
		.hps_0_h2f_axi_master_arprot                                 (hps_0_h2f_axi_master_arprot),                                                   //                                                  .arprot
		.hps_0_h2f_axi_master_arvalid                                (hps_0_h2f_axi_master_arvalid),                                                  //                                                  .arvalid
		.hps_0_h2f_axi_master_arready                                (hps_0_h2f_axi_master_arready),                                                  //                                                  .arready
		.hps_0_h2f_axi_master_rid                                    (hps_0_h2f_axi_master_rid),                                                      //                                                  .rid
		.hps_0_h2f_axi_master_rdata                                  (hps_0_h2f_axi_master_rdata),                                                    //                                                  .rdata
		.hps_0_h2f_axi_master_rresp                                  (hps_0_h2f_axi_master_rresp),                                                    //                                                  .rresp
		.hps_0_h2f_axi_master_rlast                                  (hps_0_h2f_axi_master_rlast),                                                    //                                                  .rlast
		.hps_0_h2f_axi_master_rvalid                                 (hps_0_h2f_axi_master_rvalid),                                                   //                                                  .rvalid
		.hps_0_h2f_axi_master_rready                                 (hps_0_h2f_axi_master_rready),                                                   //                                                  .rready
		.clk_0_clk_clk                                               (clk_clk),                                                                       //                                         clk_0_clk.clk
		.parallel_port_out_axi_reset_reset_bridge_in_reset_reset     (rst_controller_reset_out_reset),                                                // parallel_port_out_axi_reset_reset_bridge_in_reset.reset
		.parallel_port_in_axi_avalon_parallel_port_slave_address     (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_address),     //   parallel_port_in_axi_avalon_parallel_port_slave.address
		.parallel_port_in_axi_avalon_parallel_port_slave_write       (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_write),       //                                                  .write
		.parallel_port_in_axi_avalon_parallel_port_slave_read        (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_read),        //                                                  .read
		.parallel_port_in_axi_avalon_parallel_port_slave_readdata    (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_readdata),    //                                                  .readdata
		.parallel_port_in_axi_avalon_parallel_port_slave_writedata   (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_writedata),   //                                                  .writedata
		.parallel_port_in_axi_avalon_parallel_port_slave_byteenable  (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_byteenable),  //                                                  .byteenable
		.parallel_port_in_axi_avalon_parallel_port_slave_chipselect  (mm_interconnect_0_parallel_port_in_axi_avalon_parallel_port_slave_chipselect),  //                                                  .chipselect
		.parallel_port_out_axi_avalon_parallel_port_slave_address    (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_address),    //  parallel_port_out_axi_avalon_parallel_port_slave.address
		.parallel_port_out_axi_avalon_parallel_port_slave_write      (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_write),      //                                                  .write
		.parallel_port_out_axi_avalon_parallel_port_slave_read       (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_read),       //                                                  .read
		.parallel_port_out_axi_avalon_parallel_port_slave_readdata   (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_readdata),   //                                                  .readdata
		.parallel_port_out_axi_avalon_parallel_port_slave_writedata  (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_writedata),  //                                                  .writedata
		.parallel_port_out_axi_avalon_parallel_port_slave_byteenable (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_byteenable), //                                                  .byteenable
		.parallel_port_out_axi_avalon_parallel_port_slave_chipselect (mm_interconnect_0_parallel_port_out_axi_avalon_parallel_port_slave_chipselect)  //                                                  .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
